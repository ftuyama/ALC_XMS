library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.NUMERIC_STD.all;

ENTITY hp_ex01_SYNC IS
  PORT (
    INPUT  : IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
    RESET  : IN  STD_LOGIC;
    CLOCK  : IN  STD_LOGIC
  );
END ENTITY hp_ex01_SYNC;

ARCHITECTURE ALC_XMS OF hp_ex01_SYNC IS

COMPONENT hp_ex01_SYNC_Block IS
  PORT (
    INPUT  : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
  );
END COMPONENT;

  SIGNAL SSTATE : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL SOUT   : STD_LOGIC_VECTOR(5 DOWNTO 0);

BEGIN
B: hp_ex01_SYNC_Block    PORT MAP(INPUT & SSTATE, SOUT);
 
  PROCESS(CLOCK)
  BEGIN
    IF (RISING_EDGE(CLOCK)) THEN
    	SSTATE <= SOUT(5 DOWNTO 5);
    	OUTPUT <= SOUT(4 DOWNTO 0);
    END IF;
  END PROCESS;
END ALC_XMS;
