library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.NUMERIC_STD.all;

ENTITY pe_rcv_ifc_SYNC IS
  PORT (
    INPUT  : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    RESET  : IN  STD_LOGIC;
    CLOCK  : IN  STD_LOGIC
  );
END ENTITY pe_rcv_ifc_SYNC;

ARCHITECTURE ALC_XMS OF pe_rcv_ifc_SYNC IS

COMPONENT pe_rcv_ifc_SYNC_Block IS
  PORT (
    INPUT  : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(10 DOWNTO 0)
  );
END COMPONENT;

  SIGNAL SSTATE : STD_LOGIC_VECTOR(6 DOWNTO 0);
  SIGNAL SOUT   : STD_LOGIC_VECTOR(10 DOWNTO 0);

BEGIN
B: pe_rcv_ifc_SYNC_Block    PORT MAP(INPUT & SSTATE, SOUT);
 
  PROCESS(CLOCK)
  BEGIN
    IF (RISING_EDGE(CLOCK)) THEN
    	SSTATE <= SOUT(10 DOWNTO 4);
    	OUTPUT <= SOUT(3 DOWNTO 0);
    END IF;
  END PROCESS;
END ALC_XMS;
