library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.NUMERIC_STD.all;

ENTITY sc_control IS
  PORT (
    INPUT  : IN  STD_LOGIC_VECTOR(12 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(16 DOWNTO 0);
    STATE  : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
    RSTATE : IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
    RESET  : IN  STD_LOGIC;
    IN_DELAY  : IN  STD_LOGIC;
    OUT_DELAY : OUT STD_LOGIC
  );
END ENTITY sc_control;

ARCHITECTURE ALC_XMS OF sc_control IS

COMPONENT FGC_Block IS
  PORT (
    INPUT  : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC
  );
END COMPONENT;

COMPONENT NSTATE_Block IS
  PORT (
    INPUT  : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
  );
END COMPONENT;

COMPONENT OUT_Block IS
  PORT (
    INPUT  : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(16 DOWNTO 0)
  );
END COMPONENT;

COMPONENT D_Latch IS
  Port (
    EN : in  STD_LOGIC;
    D  : in  STD_LOGIC;
    Q  : out STD_LOGIC
  );
END COMPONENT;

  SIGNAL SSTATE : STD_LOGIC_VECTOR(4 DOWNTO 0);
  SIGNAL SNSTATE: STD_LOGIC_VECTOR(4 DOWNTO 0);
  SIGNAL SLSTATE: STD_LOGIC_VECTOR(4 DOWNTO 0);
  SIGNAL SSOUT  : STD_LOGIC_VECTOR(16 DOWNTO 0);
  SIGNAL SOUT   : STD_LOGIC_VECTOR(16 DOWNTO 0);

BEGIN
B1: FGC_Block    PORT MAP(INPUT & SSTATE, OUT_DELAY);
B2: NSTATE_Block PORT MAP(INPUT & SSTATE, SNSTATE);
B3: OUT_Block    PORT MAP(INPUT & SSTATE, SOUT);
STT0: D_Latch    PORT MAP(IN_DELAY OR RESET, SLSTATE(0), SSTATE(0));
STT1: D_Latch    PORT MAP(IN_DELAY OR RESET, SLSTATE(1), SSTATE(1));
STT2: D_Latch    PORT MAP(IN_DELAY OR RESET, SLSTATE(2), SSTATE(2));
STT3: D_Latch    PORT MAP(IN_DELAY OR RESET, SLSTATE(3), SSTATE(3));
STT4: D_Latch    PORT MAP(IN_DELAY OR RESET, SLSTATE(4), SSTATE(4));
OUT0: D_Latch    PORT MAP(SSOUT(0) XOR SOUT(0), SOUT(0), OUTPUT(0));
OUT1: D_Latch    PORT MAP(SSOUT(1) XOR SOUT(1), SOUT(1), OUTPUT(1));
OUT2: D_Latch    PORT MAP(SSOUT(2) XOR SOUT(2), SOUT(2), OUTPUT(2));
OUT3: D_Latch    PORT MAP(SSOUT(3) XOR SOUT(3), SOUT(3), OUTPUT(3));
OUT4: D_Latch    PORT MAP(SSOUT(4) XOR SOUT(4), SOUT(4), OUTPUT(4));
OUT5: D_Latch    PORT MAP(SSOUT(5) XOR SOUT(5), SOUT(5), OUTPUT(5));
OUT6: D_Latch    PORT MAP(SSOUT(6) XOR SOUT(6), SOUT(6), OUTPUT(6));
OUT7: D_Latch    PORT MAP(SSOUT(7) XOR SOUT(7), SOUT(7), OUTPUT(7));
OUT8: D_Latch    PORT MAP(SSOUT(8) XOR SOUT(8), SOUT(8), OUTPUT(8));
OUT9: D_Latch    PORT MAP(SSOUT(9) XOR SOUT(9), SOUT(9), OUTPUT(9));
OUT10: D_Latch    PORT MAP(SSOUT(10) XOR SOUT(10), SOUT(10), OUTPUT(10));
OUT11: D_Latch    PORT MAP(SSOUT(11) XOR SOUT(11), SOUT(11), OUTPUT(11));
OUT12: D_Latch    PORT MAP(SSOUT(12) XOR SOUT(12), SOUT(12), OUTPUT(12));
OUT13: D_Latch    PORT MAP(SSOUT(13) XOR SOUT(13), SOUT(13), OUTPUT(13));
OUT14: D_Latch    PORT MAP(SSOUT(14) XOR SOUT(14), SOUT(14), OUTPUT(14));
OUT15: D_Latch    PORT MAP(SSOUT(15) XOR SOUT(15), SOUT(15), OUTPUT(15));
OUT16: D_Latch    PORT MAP(SSOUT(16) XOR SOUT(16), SOUT(16), OUTPUT(16));
 
  PROCESS(INPUT, RSTATE, RESET, IN_DELAY)
  BEGIN
    OUTPUT <= SSOUT;
    IF (RESET = '1') THEN
      SLSTATE <= RSTATE;
    ELSE
      SLSTATE <= SNSTATE;
    END IF;
    STATE <= SSTATE;
  END PROCESS;
END ALC_XMS;
