library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.NUMERIC_STD.all;

ENTITY pscsi_SYNC_Block IS
  PORT (
    INPUT : IN  STD_LOGIC_VECTOR(17 DOWNTO 0);
    OUTPUT: OUT STD_LOGIC_VECTOR(12 DOWNTO 0)
  );
END pscsi_SYNC_Block;

ARCHITECTURE version OF pscsi_SYNC_Block IS
BEGIN
  PROCESS(INPUT)
  BEGIN
     if std_match(INPUT, "010-11-1110-0-0--0") then OUTPUT <= "---------1-1-";
     elsif std_match(INPUT, "-----101--0-00000-") then OUTPUT <= "-1-------1---";
     elsif std_match(INPUT, "1--------000000-00") then OUTPUT <= "-----1-------";
     elsif std_match(INPUT, "----1-0----0-00000") then OUTPUT <= "1------------";
     elsif std_match(INPUT, "---------00-000000") then OUTPUT <= "-1-----------";
     elsif std_match(INPUT, "------0---0-000000") then OUTPUT <= "-1-------1---";
     elsif std_match(INPUT, "----110---000-00-0") then OUTPUT <= "---1-----1-1-";
     elsif std_match(INPUT, "01-------100000--0") then OUTPUT <= "-----1---1-1-";
     elsif std_match(INPUT, "0--------000-00000") then OUTPUT <= "--1-------11-";
     elsif std_match(INPUT, "-00---1---000----0") then OUTPUT <= "---------1---";
     elsif std_match(INPUT, "-0----1---000-00-0") then OUTPUT <= "---1-------1-";
     elsif std_match(INPUT, "0-0-11-11--1------") then OUTPUT <= "-1-------11--";
     elsif std_match(INPUT, "0---0-----00-0000-") then OUTPUT <= "--1-------11-";
     elsif std_match(INPUT, "1-0-11-11-----1---") then OUTPUT <= "----1----1-1-";
     elsif std_match(INPUT, "0--------0-000-000") then OUTPUT <= "1---------11-";
     elsif std_match(INPUT, "1--------0-00000-0") then OUTPUT <= "1---------11-";
     elsif std_match(INPUT, "----0-1-----00000-") then OUTPUT <= "--1-------11-";
     elsif std_match(INPUT, "1---11-11---1-----") then OUTPUT <= "--1--------1-";
     elsif std_match(INPUT, "1--------00-0-0-00") then OUTPUT <= "----------111";
     elsif std_match(INPUT, "--00--1-111-------") then OUTPUT <= "1-------1-11-";
     elsif std_match(INPUT, "-1--11---1---1----") then OUTPUT <= "------1----1-";
     elsif std_match(INPUT, "1----1-1-1-1------") then OUTPUT <= "--1--------1-";
     elsif std_match(INPUT, "01--1----1--1-----") then OUTPUT <= "----1------1-";
     elsif std_match(INPUT, "01--11----------1-") then OUTPUT <= "-----1---1-1-";
     elsif std_match(INPUT, "0-0-11---------1--") then OUTPUT <= "-----1---1-1-";
     elsif std_match(INPUT, "1------110-------1") then OUTPUT <= "-------1-1-1-";
     elsif std_match(INPUT, "01---0---------00-") then OUTPUT <= "---1------11-";
     elsif std_match(INPUT, "-0---01----1------") then OUTPUT <= "-------1---1-";
     elsif std_match(INPUT, "1---1----1------1-") then OUTPUT <= "------1----1-";
     elsif std_match(INPUT, "----0-0----00-----") then OUTPUT <= "1----------1-";
     elsif std_match(INPUT, "0-----1--1----1---") then OUTPUT <= "----1------1-";
     elsif std_match(INPUT, "0-----10-1--------") then OUTPUT <= "-------1---1-";
     elsif std_match(INPUT, "----110-------1---") then OUTPUT <= "----1----1-1-";
     elsif std_match(INPUT, "1--------1----1---") then OUTPUT <= "----------1--";
     elsif std_match(INPUT, "-01-------1-------") then OUTPUT <= "----1------1-";
     elsif std_match(INPUT, "1-------11-----1--") then OUTPUT <= "1-------1-11-";
     elsif std_match(INPUT, "0-----1-01--------") then OUTPUT <= "1---------11-";
     elsif std_match(INPUT, "-0----1--------1--") then OUTPUT <= "-----1-----1-";
     elsif std_match(INPUT, "-----00----0------") then OUTPUT <= "-------1---1-";
     elsif std_match(INPUT, "-0----1-----1-----") then OUTPUT <= "--1--------1-";
     elsif std_match(INPUT, "0------0---------1") then OUTPUT <= "-------1---1-";
     elsif std_match(INPUT, "------1--1-------1") then OUTPUT <= "-------1---1-";
     elsif std_match(INPUT, "0------1-0-------1") then OUTPUT <= "-1-------111-";
     elsif std_match(INPUT, "1--------1--1-----") then OUTPUT <= "--1--------1-";
     elsif std_match(INPUT, "----0---------1---") then OUTPUT <= "----------1--";
     elsif std_match(INPUT, "011---------------") then OUTPUT <= "-1--------11-";
     elsif std_match(INPUT, "--------00--1-----") then OUTPUT <= "-----1----111";
     elsif std_match(INPUT, "-------0-0--1-----") then OUTPUT <= "-1--------111";
     elsif std_match(INPUT, "0----0---0--------") then OUTPUT <= "---1------11-";
     elsif std_match(INPUT, "-----0---0--1-----") then OUTPUT <= "-1--------111";
     elsif std_match(INPUT, "0---0----0--------") then OUTPUT <= "--1-------11-";
     elsif std_match(INPUT, "0--------0-1------") then OUTPUT <= "---------111-";
     elsif std_match(INPUT, "1-------0---0-----") then OUTPUT <= "-----1----111";
     elsif std_match(INPUT, "1---0----0--------") then OUTPUT <= "---1------111";
     elsif std_match(INPUT, "1------0----0-----") then OUTPUT <= "-1--------111";
     elsif std_match(INPUT, "1---0-------0-----") then OUTPUT <= "---1------111";
     elsif std_match(INPUT, "1----0------0-----") then OUTPUT <= "-1--------111";
     elsif std_match(INPUT, "-0----------------") then OUTPUT <= "----------1--";
     elsif std_match(INPUT, "---------0---1----") then OUTPUT <= "---1------11-";
     elsif std_match(INPUT, "1-1---------------") then OUTPUT <= "----1-----11-";
     elsif std_match(INPUT, "---1--------------") then OUTPUT <= "-------1--11-";
     elsif std_match(INPUT, "000001011110000000") then OUTPUT <= "-000000000--0";
     elsif std_match(INPUT, "000001011101000000") then OUTPUT <= "0-0000000--00";
     elsif std_match(INPUT, "000001011100100000") then OUTPUT <= "00-0000000--0";
     elsif std_match(INPUT, "000001011100010000") then OUTPUT <= "-000000000--0";
     elsif std_match(INPUT, "000001011100001000") then OUTPUT <= "-000000000--0";
     elsif std_match(INPUT, "000001011100000100") then OUTPUT <= "-000000000--0";
     elsif std_match(INPUT, "000001011100000010") then OUTPUT <= "-000000000--0";
     elsif std_match(INPUT, "000001111101000000") then OUTPUT <= "00-0000000--0";
     elsif std_match(INPUT, "000001111100100000") then OUTPUT <= "00-0000000--0";
     elsif std_match(INPUT, "000001111100010000") then OUTPUT <= "000-00000---0";
     elsif std_match(INPUT, "000001111100001000") then OUTPUT <= "0000-0000---0";
     elsif std_match(INPUT, "000001111100000100") then OUTPUT <= "00000-000---0";
     elsif std_match(INPUT, "000001111100000010") then OUTPUT <= "000-00000---0";
     elsif std_match(INPUT, "000010011100000001") then OUTPUT <= "0000000-00--0";
     elsif std_match(INPUT, "000010011101000000") then OUTPUT <= "0-0000000--00";
     elsif std_match(INPUT, "000010011100010000") then OUTPUT <= "0000000-00--0";
     elsif std_match(INPUT, "000010011100001000") then OUTPUT <= "0000000-00--0";
     elsif std_match(INPUT, "000010011100000100") then OUTPUT <= "0000000-00--0";
     elsif std_match(INPUT, "000010011100000010") then OUTPUT <= "0000000-00--0";
     elsif std_match(INPUT, "000010111100000001") then OUTPUT <= "0000000-00--0";
     elsif std_match(INPUT, "000010111101000000") then OUTPUT <= "0000000-00--0";
     elsif std_match(INPUT, "000010111100010000") then OUTPUT <= "000-00000---0";
     elsif std_match(INPUT, "000010111100001000") then OUTPUT <= "0000-0000---0";
     elsif std_match(INPUT, "000010111100000100") then OUTPUT <= "00000-000---0";
     elsif std_match(INPUT, "000010111100000010") then OUTPUT <= "000-00000---0";
     elsif std_match(INPUT, "000011001100000001") then OUTPUT <= "0000000-00--0";
     elsif std_match(INPUT, "000011001101000000") then OUTPUT <= "0-0000000--00";
     elsif std_match(INPUT, "000011010101000000") then OUTPUT <= "0-0000000--00";
     elsif std_match(INPUT, "000011011110000000") then OUTPUT <= "-000000000-00";
     elsif std_match(INPUT, "000011011100000001") then OUTPUT <= "0-0000000--00";
     elsif std_match(INPUT, "000011011101000000") then OUTPUT <= "0-0000000--00";
     elsif std_match(INPUT, "000011011100100000") then OUTPUT <= "-000000000-00";
     elsif std_match(INPUT, "000011011100010000") then OUTPUT <= "000-00000---0";
     elsif std_match(INPUT, "000011011100001000") then OUTPUT <= "0000-0000---0";
     elsif std_match(INPUT, "000011011100000100") then OUTPUT <= "00000-000---0";
     elsif std_match(INPUT, "000011011100000010") then OUTPUT <= "000-00000---0";
     elsif std_match(INPUT, "000011101100000001") then OUTPUT <= "0000000-00--0";
     elsif std_match(INPUT, "000011101101000000") then OUTPUT <= "0000000-00--0";
     elsif std_match(INPUT, "000011110110000000") then OUTPUT <= "-000000000--0";
     elsif std_match(INPUT, "000011110101000000") then OUTPUT <= "-000000000--0";
     elsif std_match(INPUT, "000011111110000000") then OUTPUT <= "-0000000-0--0";
     elsif std_match(INPUT, "000011111100000001") then OUTPUT <= "0000000-00--0";
     elsif std_match(INPUT, "000011111101000000") then OUTPUT <= "0-0000000--00";
     elsif std_match(INPUT, "000011111100100000") then OUTPUT <= "00-0000000--0";
     elsif std_match(INPUT, "000011111100010000") then OUTPUT <= "000-00000---0";
     elsif std_match(INPUT, "000011111100001000") then OUTPUT <= "0000-0000---0";
     elsif std_match(INPUT, "000011111100000100") then OUTPUT <= "00000-000---0";
     elsif std_match(INPUT, "000011111100000010") then OUTPUT <= "000-00000---0";
     elsif std_match(INPUT, "000111111110000000") then OUTPUT <= "0000000-00--0";
     elsif std_match(INPUT, "000111111100000001") then OUTPUT <= "0000000-00--0";
     elsif std_match(INPUT, "001011111110000000") then OUTPUT <= "0000-00000--0";
     elsif std_match(INPUT, "001011111100010000") then OUTPUT <= "000-000000--0";
     elsif std_match(INPUT, "001011111100001000") then OUTPUT <= "0000-00000--0";
     elsif std_match(INPUT, "001011111100000100") then OUTPUT <= "00000-0000--0";
     elsif std_match(INPUT, "001011111100000010") then OUTPUT <= "000-000000--0";
     elsif std_match(INPUT, "010001111000100000") then OUTPUT <= "00-0000000--0";
     elsif std_match(INPUT, "010001111000000100") then OUTPUT <= "00-0000000--0";
     elsif std_match(INPUT, "010001111000000010") then OUTPUT <= "00-0000000--0";
     elsif std_match(INPUT, "010001111101000000") then OUTPUT <= "00-0000000--0";
     elsif std_match(INPUT, "010001111100100000") then OUTPUT <= "00-0000000--0";
     elsif std_match(INPUT, "010001111100001000") then OUTPUT <= "0000-00000--0";
     elsif std_match(INPUT, "010001111100000100") then OUTPUT <= "00000-000-0-0";
     elsif std_match(INPUT, "010001111100000010") then OUTPUT <= "00000-000-0-0";
     elsif std_match(INPUT, "010010111000010000") then OUTPUT <= "000-000000--0";
     elsif std_match(INPUT, "010010111000000100") then OUTPUT <= "000-000000--0";
     elsif std_match(INPUT, "010010111000000010") then OUTPUT <= "000-000000--0";
     elsif std_match(INPUT, "010010111101000000") then OUTPUT <= "000-000000--0";
     elsif std_match(INPUT, "010010111100010000") then OUTPUT <= "000-000000--0";
     elsif std_match(INPUT, "010010111100000100") then OUTPUT <= "00000-000-0-0";
     elsif std_match(INPUT, "010010111100000010") then OUTPUT <= "00000-000-0-0";
     elsif std_match(INPUT, "010011101000000001") then OUTPUT <= "0000000-000-0";
     elsif std_match(INPUT, "010011101001000000") then OUTPUT <= "0-0000000---0";
     elsif std_match(INPUT, "010011101100000001") then OUTPUT <= "0000000-000-0";
     elsif std_match(INPUT, "010011101101000000") then OUTPUT <= "0000000-000-0";
     elsif std_match(INPUT, "010011110001000000") then OUTPUT <= "0-0000000---0";
     elsif std_match(INPUT, "010011110110000000") then OUTPUT <= "-000000000--0";
     elsif std_match(INPUT, "010011110101000000") then OUTPUT <= "-000000000--0";
     elsif std_match(INPUT, "010011111010000000") then OUTPUT <= "-000000000--0";
     elsif std_match(INPUT, "010011111000000001") then OUTPUT <= "0-0000000---0";
     elsif std_match(INPUT, "010011111001000000") then OUTPUT <= "0-0000000---0";
     elsif std_match(INPUT, "010011111000100000") then OUTPUT <= "00-0000000--0";
     elsif std_match(INPUT, "010011111000010000") then OUTPUT <= "000-000000--0";
     elsif std_match(INPUT, "010011111000001000") then OUTPUT <= "-000000000--0";
     elsif std_match(INPUT, "010011111000000100") then OUTPUT <= "00000-000-0-0";
     elsif std_match(INPUT, "010011111000000010") then OUTPUT <= "00000-000-0-0";
     elsif std_match(INPUT, "010011111110000000") then OUTPUT <= "-0000000-0--0";
     elsif std_match(INPUT, "010011111100000001") then OUTPUT <= "0000000-000-0";
     elsif std_match(INPUT, "010011111101000000") then OUTPUT <= "0-0000000---0";
     elsif std_match(INPUT, "010011111100100000") then OUTPUT <= "0000-000000-0";
     elsif std_match(INPUT, "010011111100010000") then OUTPUT <= "000000-00-0-0";
     elsif std_match(INPUT, "010011111100001000") then OUTPUT <= "0000-000000-0";
     elsif std_match(INPUT, "010011111100000100") then OUTPUT <= "00000-000-0-0";
     elsif std_match(INPUT, "010011111100000010") then OUTPUT <= "00000-000-0-0";
     elsif std_match(INPUT, "010111111110000000") then OUTPUT <= "0000000-00--0";
     elsif std_match(INPUT, "010111111100000001") then OUTPUT <= "0000000-00--0";
     elsif std_match(INPUT, "011011111110000000") then OUTPUT <= "0-00000000--0";
     elsif std_match(INPUT, "011011111101000000") then OUTPUT <= "0-00000000--0";
     elsif std_match(INPUT, "110001111000100000") then OUTPUT <= "000-000000---";
     elsif std_match(INPUT, "110001111000010000") then OUTPUT <= "000-000000---";
     elsif std_match(INPUT, "110001111100100000") then OUTPUT <= "00-00000000-0";
     elsif std_match(INPUT, "110001111100010000") then OUTPUT <= "000-000000---";
     elsif std_match(INPUT, "110001111100001000") then OUTPUT <= "000-000000---";
     elsif std_match(INPUT, "110001111100000010") then OUTPUT <= "000-000000---";
     elsif std_match(INPUT, "110010111001000000") then OUTPUT <= "0-00000000---";
     elsif std_match(INPUT, "110010111000100000") then OUTPUT <= "0-00000000---";
     elsif std_match(INPUT, "110010111101000000") then OUTPUT <= "0-00000000---";
     elsif std_match(INPUT, "110010111100100000") then OUTPUT <= "00-00000000-0";
     elsif std_match(INPUT, "110010111100001000") then OUTPUT <= "0-00000000---";
     elsif std_match(INPUT, "110011101000000001") then OUTPUT <= "0-00000000---";
     elsif std_match(INPUT, "110011101001000000") then OUTPUT <= "0-00000000---";
     elsif std_match(INPUT, "110011101000100000") then OUTPUT <= "0-00000000---";
     elsif std_match(INPUT, "110011101000001000") then OUTPUT <= "0-00000000---";
     elsif std_match(INPUT, "110011101101000000") then OUTPUT <= "0-00000000---";
     elsif std_match(INPUT, "110011101100100000") then OUTPUT <= "00-00000000-0";
     elsif std_match(INPUT, "110011110000000001") then OUTPUT <= "00000-0000---";
     elsif std_match(INPUT, "110011110000100000") then OUTPUT <= "00000-0000---";
     elsif std_match(INPUT, "110011110000001000") then OUTPUT <= "00000-0000---";
     elsif std_match(INPUT, "110011110000000100") then OUTPUT <= "00000-0000---";
     elsif std_match(INPUT, "110011110100100000") then OUTPUT <= "00-00000000-0";
     elsif std_match(INPUT, "110011110100000100") then OUTPUT <= "00000-0000---";
     elsif std_match(INPUT, "110011111010000000") then OUTPUT <= "-000000000--0";
     elsif std_match(INPUT, "110011111000000001") then OUTPUT <= "0000000-0-0-0";
     elsif std_match(INPUT, "110011111001000000") then OUTPUT <= "0-00000000---";
     elsif std_match(INPUT, "110011111000100000") then OUTPUT <= "00-00000000-0";
     elsif std_match(INPUT, "110011111000010000") then OUTPUT <= "000-000000---";
     elsif std_match(INPUT, "110011111000001000") then OUTPUT <= "0000-0000-0-0";
     elsif std_match(INPUT, "110011111000000100") then OUTPUT <= "00000-0000---";
     elsif std_match(INPUT, "110011111000000010") then OUTPUT <= "-000000000--0";
     elsif std_match(INPUT, "110011111110000000") then OUTPUT <= "-0000000-0--0";
     elsif std_match(INPUT, "110011111100000001") then OUTPUT <= "0000000-000-0";
     elsif std_match(INPUT, "110011111101000000") then OUTPUT <= "00-00000000-0";
     elsif std_match(INPUT, "110011111100100000") then OUTPUT <= "00-00000000-0";
     elsif std_match(INPUT, "110011111100010000") then OUTPUT <= "000000-0000-0";
     elsif std_match(INPUT, "110011111100001000") then OUTPUT <= "0000-0000---0";
     elsif std_match(INPUT, "110011111100000100") then OUTPUT <= "-0000000-0--0";
     elsif std_match(INPUT, "110011111100000010") then OUTPUT <= "000000-0000-0";
     elsif std_match(INPUT, "110111111110000000") then OUTPUT <= "0000000-00--0";
     elsif std_match(INPUT, "110111111100000001") then OUTPUT <= "0000000-00--0";
     elsif std_match(INPUT, "111011111110000000") then OUTPUT <= "0000-00000--0";
     elsif std_match(INPUT, "111011111100001000") then OUTPUT <= "0000-00000--0";
     else OUTPUT <= "-------------";
    END if;

  END PROCESS;
END version;
