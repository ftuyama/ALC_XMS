library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.NUMERIC_STD.all;

ENTITY call_proc_SYNC IS
  PORT (
    INPUT  : IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
    RESET  : IN  STD_LOGIC;
    CLOCK  : IN  STD_LOGIC
  );
END ENTITY call_proc_SYNC;

ARCHITECTURE ALC_XMS OF call_proc_SYNC IS

COMPONENT call_proc_SYNC_Block IS
  PORT (
    INPUT  : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
  );
END COMPONENT;

  SIGNAL SSTATE : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL SOUT   : STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN
B: call_proc_SYNC_Block    PORT MAP(INPUT & SSTATE, SOUT);
 
  PROCESS(CLOCK)
  BEGIN
    IF (RISING_EDGE(CLOCK)) THEN
    	SSTATE <= SOUT(3 DOWNTO 3);
    	OUTPUT <= SOUT(2 DOWNTO 0);
    END IF;
  END PROCESS;
END ALC_XMS;
