library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.NUMERIC_STD.all;

ENTITY hp_ex01_SYNC IS
  PORT (
    INPUT  : IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
    RESET  : IN  STD_LOGIC
  );
END ENTITY hp_ex01_SYNC;

ARCHITECTURE ALC_XMS OF hp_ex01_SYNC IS

COMPONENT hp_ex01_SYNC_Block IS
  PORT (
    INPUT  : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
  );
END COMPONENT;

COMPONENT D_Latch IS
  Port (
    EN : in  STD_LOGIC;
    D  : in  STD_LOGIC;
    Q  : out STD_LOGIC
  );
END COMPONENT;

  SIGNAL SSTATE : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL SOUT   : STD_LOGIC_VECTOR(5 DOWNTO 0);
  SIGNAL HIGH	 : STD_LOGIC;
BEGIN
B: hp_ex01_SYNC_Block    PORT MAP(INPUT & SSTATE, SOUT);
STT0: D_Latch    PORT MAP(RESET, SOUT(0), HIGH);
OUT1: D_Latch    PORT MAP(RESET, SOUT(1), HIGH);
OUT2: D_Latch    PORT MAP(RESET, SOUT(2), HIGH);
OUT3: D_Latch    PORT MAP(RESET, SOUT(3), HIGH);
OUT4: D_Latch    PORT MAP(RESET, SOUT(4), HIGH);
OUT5: D_Latch    PORT MAP(RESET, SOUT(5), HIGH);
 
  PROCESS(INPUT)
  BEGIN
  	 HIGH <= '1';
    SSTATE <= SOUT(5 DOWNTO 5);
    OUTPUT <= SOUT(4 DOWNTO 0);
  END PROCESS;
END ALC_XMS;
