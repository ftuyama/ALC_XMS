library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.NUMERIC_STD.all;

ENTITY re_setup_SYNC IS
  PORT (
    INPUT  : IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    RESET  : IN  STD_LOGIC
  );
END ENTITY re_setup_SYNC;

ARCHITECTURE ALC_XMS OF re_setup_SYNC IS

COMPONENT re_setup_SYNC_Block IS
  PORT (
    INPUT  : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
  );
END COMPONENT;

COMPONENT D_Latch IS
  Port (
    EN : in  STD_LOGIC;
    D  : in  STD_LOGIC;
    Q  : out STD_LOGIC
  );
END COMPONENT;

  SIGNAL SSTATE : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL SOUT   : STD_LOGIC_VECTOR(2 DOWNTO 0);
  SIGNAL HIGH	 : STD_LOGIC;
BEGIN
B: re_setup_SYNC_Block    PORT MAP(INPUT & SSTATE, SOUT);
STT0: D_Latch    PORT MAP(RESET, SOUT(0), HIGH);
OUT1: D_Latch    PORT MAP(RESET, SOUT(1), HIGH);
OUT2: D_Latch    PORT MAP(RESET, SOUT(2), HIGH);
 
  PROCESS(INPUT)
  BEGIN
  	 HIGH <= '1';
    SSTATE <= SOUT(2 DOWNTO 2);
    OUTPUT <= SOUT(1 DOWNTO 0);
  END PROCESS;
END ALC_XMS;
