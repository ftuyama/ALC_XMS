library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.NUMERIC_STD.all;

ENTITY OUT_Block IS
  PORT (
    INPUT : IN  STD_LOGIC_VECTOR(17 DOWNTO 0);
    OUTPUT: OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
  );
END OUT_Block;

ARCHITECTURE version OF OUT_Block IS
BEGIN
  PROCESS(INPUT)
  BEGIN
     if std_match(INPUT, "000001011110000000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000001011101000000") then OUTPUT <= "01100";
     elsif std_match(INPUT, "000001011100100000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000001011100010000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000001011100001000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000001011100000100") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000001011100000010") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000001111101000000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000001111100100000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000001111100010000") then OUTPUT <= "01110";
     elsif std_match(INPUT, "000001111100001000") then OUTPUT <= "01110";
     elsif std_match(INPUT, "000001111100000100") then OUTPUT <= "01110";
     elsif std_match(INPUT, "000001111100000010") then OUTPUT <= "01110";
     elsif std_match(INPUT, "000010011100000001") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000010011101000000") then OUTPUT <= "01100";
     elsif std_match(INPUT, "000010011100010000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000010011100001000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000010011100000100") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000010011100000010") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000010111100000001") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000010111101000000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000010111100010000") then OUTPUT <= "01110";
     elsif std_match(INPUT, "000010111100001000") then OUTPUT <= "01110";
     elsif std_match(INPUT, "000010111100000100") then OUTPUT <= "01110";
     elsif std_match(INPUT, "000010111100000010") then OUTPUT <= "01110";
     elsif std_match(INPUT, "000011001100000001") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000011001101000000") then OUTPUT <= "01100";
     elsif std_match(INPUT, "000011010101000000") then OUTPUT <= "01100";
     elsif std_match(INPUT, "000011011110000000") then OUTPUT <= "00100";
     elsif std_match(INPUT, "000011011100000001") then OUTPUT <= "01100";
     elsif std_match(INPUT, "000011011101000000") then OUTPUT <= "01100";
     elsif std_match(INPUT, "000011011100100000") then OUTPUT <= "00100";
     elsif std_match(INPUT, "000011011100010000") then OUTPUT <= "01110";
     elsif std_match(INPUT, "000011011100001000") then OUTPUT <= "01110";
     elsif std_match(INPUT, "000011011100000100") then OUTPUT <= "01110";
     elsif std_match(INPUT, "000011011100000010") then OUTPUT <= "01110";
     elsif std_match(INPUT, "000011101100000001") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000011101101000000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000011110110000000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000011110101000000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000011111110000000") then OUTPUT <= "10110";
     elsif std_match(INPUT, "000011111100000001") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000011111101000000") then OUTPUT <= "01100";
     elsif std_match(INPUT, "000011111100100000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000011111100010000") then OUTPUT <= "01110";
     elsif std_match(INPUT, "000011111100001000") then OUTPUT <= "01110";
     elsif std_match(INPUT, "000011111100000100") then OUTPUT <= "01110";
     elsif std_match(INPUT, "000011111100000010") then OUTPUT <= "01110";
     elsif std_match(INPUT, "000111111110000000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "000111111100000001") then OUTPUT <= "00110";
     elsif std_match(INPUT, "001011111110000000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "001011111100010000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "001011111100001000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "001011111100000100") then OUTPUT <= "00110";
     elsif std_match(INPUT, "001011111100000010") then OUTPUT <= "00110";
     elsif std_match(INPUT, "010001111000100000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "010001111000000100") then OUTPUT <= "00110";
     elsif std_match(INPUT, "010001111000000010") then OUTPUT <= "00110";
     elsif std_match(INPUT, "010001111101000000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "010001111100100000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "010001111100001000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "010001111100000100") then OUTPUT <= "01010";
     elsif std_match(INPUT, "010001111100000010") then OUTPUT <= "01010";
     elsif std_match(INPUT, "010010111000010000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "010010111000000100") then OUTPUT <= "00110";
     elsif std_match(INPUT, "010010111000000010") then OUTPUT <= "00110";
     elsif std_match(INPUT, "010010111101000000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "010010111100010000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "010010111100000100") then OUTPUT <= "01010";
     elsif std_match(INPUT, "010010111100000010") then OUTPUT <= "01010";
     elsif std_match(INPUT, "010011101000000001") then OUTPUT <= "00010";
     elsif std_match(INPUT, "010011101001000000") then OUTPUT <= "01110";
     elsif std_match(INPUT, "010011101100000001") then OUTPUT <= "00010";
     elsif std_match(INPUT, "010011101101000000") then OUTPUT <= "00010";
     elsif std_match(INPUT, "010011110001000000") then OUTPUT <= "01110";
     elsif std_match(INPUT, "010011110110000000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "010011110101000000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "010011111010000000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "010011111000000001") then OUTPUT <= "01110";
     elsif std_match(INPUT, "010011111001000000") then OUTPUT <= "01110";
     elsif std_match(INPUT, "010011111000100000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "010011111000010000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "010011111000001000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "010011111000000100") then OUTPUT <= "01010";
     elsif std_match(INPUT, "010011111000000010") then OUTPUT <= "01010";
     elsif std_match(INPUT, "010011111110000000") then OUTPUT <= "10110";
     elsif std_match(INPUT, "010011111100000001") then OUTPUT <= "00010";
     elsif std_match(INPUT, "010011111101000000") then OUTPUT <= "01110";
     elsif std_match(INPUT, "010011111100100000") then OUTPUT <= "00010";
     elsif std_match(INPUT, "010011111100010000") then OUTPUT <= "01010";
     elsif std_match(INPUT, "010011111100001000") then OUTPUT <= "00010";
     elsif std_match(INPUT, "010011111100000100") then OUTPUT <= "01010";
     elsif std_match(INPUT, "010011111100000010") then OUTPUT <= "01010";
     elsif std_match(INPUT, "010111111110000000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "010111111100000001") then OUTPUT <= "00110";
     elsif std_match(INPUT, "011011111110000000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "011011111101000000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "110001111000100000") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110001111000010000") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110001111100100000") then OUTPUT <= "00010";
     elsif std_match(INPUT, "110001111100010000") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110001111100001000") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110001111100000010") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110010111001000000") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110010111000100000") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110010111101000000") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110010111100100000") then OUTPUT <= "00010";
     elsif std_match(INPUT, "110010111100001000") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110011101000000001") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110011101001000000") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110011101000100000") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110011101000001000") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110011101101000000") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110011101100100000") then OUTPUT <= "00010";
     elsif std_match(INPUT, "110011110000000001") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110011110000100000") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110011110000001000") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110011110000000100") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110011110100100000") then OUTPUT <= "00010";
     elsif std_match(INPUT, "110011110100000100") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110011111010000000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "110011111000000001") then OUTPUT <= "01010";
     elsif std_match(INPUT, "110011111001000000") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110011111000100000") then OUTPUT <= "00010";
     elsif std_match(INPUT, "110011111000010000") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110011111000001000") then OUTPUT <= "01010";
     elsif std_match(INPUT, "110011111000000100") then OUTPUT <= "00111";
     elsif std_match(INPUT, "110011111000000010") then OUTPUT <= "00110";
     elsif std_match(INPUT, "110011111110000000") then OUTPUT <= "10110";
     elsif std_match(INPUT, "110011111100000001") then OUTPUT <= "00010";
     elsif std_match(INPUT, "110011111101000000") then OUTPUT <= "00010";
     elsif std_match(INPUT, "110011111100100000") then OUTPUT <= "00010";
     elsif std_match(INPUT, "110011111100010000") then OUTPUT <= "00010";
     elsif std_match(INPUT, "110011111100001000") then OUTPUT <= "01110";
     elsif std_match(INPUT, "110011111100000100") then OUTPUT <= "10110";
     elsif std_match(INPUT, "110011111100000010") then OUTPUT <= "00010";
     elsif std_match(INPUT, "110111111110000000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "110111111100000001") then OUTPUT <= "00110";
     elsif std_match(INPUT, "111011111110000000") then OUTPUT <= "00110";
     elsif std_match(INPUT, "111011111100001000") then OUTPUT <= "00110";
     else OUTPUT <= "-----";
    END if;

  END PROCESS;
END version;
