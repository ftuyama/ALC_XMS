library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.NUMERIC_STD.all;

ENTITY sc_control_SYNC IS
  PORT (
    INPUT  : IN  STD_LOGIC_VECTOR(12 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(16 DOWNTO 0);
    RESET  : IN  STD_LOGIC
  );
END ENTITY sc_control_SYNC;

ARCHITECTURE ALC_XMS OF sc_control_SYNC IS

COMPONENT sc_control_SYNC_Block IS
  PORT (
    INPUT  : IN STD_LOGIC_VECTOR(30 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(34 DOWNTO 0)
  );
END COMPONENT;

COMPONENT D_Latch IS
  Port (
    EN : in  STD_LOGIC;
    D  : in  STD_LOGIC;
    Q  : out STD_LOGIC
  );
END COMPONENT;

  SIGNAL SSTATE : STD_LOGIC_VECTOR(17 DOWNTO 0);
  SIGNAL SOUT   : STD_LOGIC_VECTOR(34 DOWNTO 0);
  SIGNAL HIGH	 : STD_LOGIC;
BEGIN
B: sc_control_SYNC_Block    PORT MAP(INPUT & SSTATE, SOUT);
STT0: D_Latch    PORT MAP(RESET, SOUT(0), HIGH);
STT1: D_Latch    PORT MAP(RESET, SOUT(1), HIGH);
STT2: D_Latch    PORT MAP(RESET, SOUT(2), HIGH);
STT3: D_Latch    PORT MAP(RESET, SOUT(3), HIGH);
STT4: D_Latch    PORT MAP(RESET, SOUT(4), HIGH);
STT5: D_Latch    PORT MAP(RESET, SOUT(5), HIGH);
STT6: D_Latch    PORT MAP(RESET, SOUT(6), HIGH);
STT7: D_Latch    PORT MAP(RESET, SOUT(7), HIGH);
STT8: D_Latch    PORT MAP(RESET, SOUT(8), HIGH);
STT9: D_Latch    PORT MAP(RESET, SOUT(9), HIGH);
STT10: D_Latch    PORT MAP(RESET, SOUT(10), HIGH);
STT11: D_Latch    PORT MAP(RESET, SOUT(11), HIGH);
STT12: D_Latch    PORT MAP(RESET, SOUT(12), HIGH);
STT13: D_Latch    PORT MAP(RESET, SOUT(13), HIGH);
STT14: D_Latch    PORT MAP(RESET, SOUT(14), HIGH);
STT15: D_Latch    PORT MAP(RESET, SOUT(15), HIGH);
STT16: D_Latch    PORT MAP(RESET, SOUT(16), HIGH);
STT17: D_Latch    PORT MAP(RESET, SOUT(17), HIGH);
OUT18: D_Latch    PORT MAP(RESET, SOUT(18), HIGH);
OUT19: D_Latch    PORT MAP(RESET, SOUT(19), HIGH);
OUT20: D_Latch    PORT MAP(RESET, SOUT(20), HIGH);
OUT21: D_Latch    PORT MAP(RESET, SOUT(21), HIGH);
OUT22: D_Latch    PORT MAP(RESET, SOUT(22), HIGH);
OUT23: D_Latch    PORT MAP(RESET, SOUT(23), HIGH);
OUT24: D_Latch    PORT MAP(RESET, SOUT(24), HIGH);
OUT25: D_Latch    PORT MAP(RESET, SOUT(25), HIGH);
OUT26: D_Latch    PORT MAP(RESET, SOUT(26), HIGH);
OUT27: D_Latch    PORT MAP(RESET, SOUT(27), HIGH);
OUT28: D_Latch    PORT MAP(RESET, SOUT(28), HIGH);
OUT29: D_Latch    PORT MAP(RESET, SOUT(29), HIGH);
OUT30: D_Latch    PORT MAP(RESET, SOUT(30), HIGH);
OUT31: D_Latch    PORT MAP(RESET, SOUT(31), HIGH);
OUT32: D_Latch    PORT MAP(RESET, SOUT(32), HIGH);
OUT33: D_Latch    PORT MAP(RESET, SOUT(33), HIGH);
OUT34: D_Latch    PORT MAP(RESET, SOUT(34), HIGH);
 
  PROCESS(INPUT)
  BEGIN
  	 HIGH <= '1';
    SSTATE <= SOUT(34 DOWNTO 17);
    OUTPUT <= SOUT(16 DOWNTO 0);
  END PROCESS;
END ALC_XMS;
