library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.NUMERIC_STD.all;

ENTITY pscsi_SYNC IS
  PORT (
    INPUT  : IN  STD_LOGIC_VECTOR(9 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
    RESET  : IN  STD_LOGIC;
    CLOCK  : IN  STD_LOGIC
  );
END ENTITY pscsi_SYNC;

ARCHITECTURE ALC_XMS OF pscsi_SYNC IS

COMPONENT pscsi_SYNC_Block IS
  PORT (
    INPUT  : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    OUTPUT : OUT STD_LOGIC_VECTOR(12 DOWNTO 0)
  );
END COMPONENT;

  SIGNAL SSTATE : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL SOUT   : STD_LOGIC_VECTOR(12 DOWNTO 0);

BEGIN
B: pscsi_SYNC_Block    PORT MAP(INPUT & SSTATE, SOUT);
 
  PROCESS(CLOCK)
  BEGIN
    IF (RISING_EDGE(CLOCK)) THEN
    	SSTATE <= SOUT(12 DOWNTO 5);
    	OUTPUT <= SOUT(4 DOWNTO 0);
    END IF;
  END PROCESS;
END ALC_XMS;
